
--tset